`include "datapath.v"

module testbench ();
  reg clk, reset;
  wire [63:0]PC, ALUResult; // Mostrar apenas as 32 bits
  wire [31:0]instruction;

  datapath Call (.clk(clk), .reset(reset), .nextPC(PC), .ALUResult(ALUResult), .instruction(instruction));

  initial begin
    $dumpfile("datapath.vcd");
    $dumpvars(0, testbench);
    $display("Exibindo os resultados:");
    $monitor("Instruction: %b\nExit PC: %b\nExit ALU: %b\n",instruction, PC, ALUResult);
  end
  initial begin
    #1; clk = 0;
    #1; clk = 1; reset = 1;
    #1; clk = 0;
    #1; clk = 1; reset = 0;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1;
    #1; clk = 0;
    #1; clk = 1; reset = 1;
    #1; clk = 0; reset = 0;
    #1;
    $finish;
  end
endmodule //

